-- soc_system_passthrough.vhd

-- Generated using ACDS version 21.1 842

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system_passthrough is
	port (
		ad1939_physical_asdata2         : in    std_logic                     := '0';             --        ad1939_physical.asdata2
		ad1939_physical_dsdata1         : out   std_logic;                                        --                       .dsdata1
		ad1939_physical_dbclk           : out   std_logic;                                        --                       .dbclk
		ad1939_physical_dlrclk          : out   std_logic;                                        --                       .dlrclk
		ad1939_physical_abclk_clk       : in    std_logic                     := '0';             --  ad1939_physical_abclk.clk
		ad1939_physical_alrclk_clk      : in    std_logic                     := '0';             -- ad1939_physical_alrclk.clk
		ad1939_physical_mclk_clk        : in    std_logic                     := '0';             --   ad1939_physical_mclk.clk
		audio_mini_leds_export          : out   std_logic_vector(3 downto 0);                     --        audio_mini_leds.export
		de10_leds_export                : out   std_logic_vector(7 downto 0);                     --              de10_leds.export
		fabric_reset_reset              : in    std_logic                     := '0';             --           fabric_reset.reset
		hps_and_fabric_reset_reset      : in    std_logic                     := '0';             --   hps_and_fabric_reset.reset
		hps_clk_clk                     : in    std_logic                     := '0';             --                hps_clk.clk
		hps_i2c0_out_data               : out   std_logic;                                        --               hps_i2c0.out_data
		hps_i2c0_sda                    : in    std_logic                     := '0';             --                       .sda
		hps_i2c0_clk_clk                : out   std_logic;                                        --           hps_i2c0_clk.clk
		hps_i2c0_scl_in_clk             : in    std_logic                     := '0';             --        hps_i2c0_scl_in.clk
		hps_io_hps_io_emac1_inst_TX_CLK : out   std_logic;                                        --                 hps_io.hps_io_emac1_inst_TX_CLK
		hps_io_hps_io_emac1_inst_TXD0   : out   std_logic;                                        --                       .hps_io_emac1_inst_TXD0
		hps_io_hps_io_emac1_inst_TXD1   : out   std_logic;                                        --                       .hps_io_emac1_inst_TXD1
		hps_io_hps_io_emac1_inst_TXD2   : out   std_logic;                                        --                       .hps_io_emac1_inst_TXD2
		hps_io_hps_io_emac1_inst_TXD3   : out   std_logic;                                        --                       .hps_io_emac1_inst_TXD3
		hps_io_hps_io_emac1_inst_RXD0   : in    std_logic                     := '0';             --                       .hps_io_emac1_inst_RXD0
		hps_io_hps_io_emac1_inst_MDIO   : inout std_logic                     := '0';             --                       .hps_io_emac1_inst_MDIO
		hps_io_hps_io_emac1_inst_MDC    : out   std_logic;                                        --                       .hps_io_emac1_inst_MDC
		hps_io_hps_io_emac1_inst_RX_CTL : in    std_logic                     := '0';             --                       .hps_io_emac1_inst_RX_CTL
		hps_io_hps_io_emac1_inst_TX_CTL : out   std_logic;                                        --                       .hps_io_emac1_inst_TX_CTL
		hps_io_hps_io_emac1_inst_RX_CLK : in    std_logic                     := '0';             --                       .hps_io_emac1_inst_RX_CLK
		hps_io_hps_io_emac1_inst_RXD1   : in    std_logic                     := '0';             --                       .hps_io_emac1_inst_RXD1
		hps_io_hps_io_emac1_inst_RXD2   : in    std_logic                     := '0';             --                       .hps_io_emac1_inst_RXD2
		hps_io_hps_io_emac1_inst_RXD3   : in    std_logic                     := '0';             --                       .hps_io_emac1_inst_RXD3
		hps_io_hps_io_sdio_inst_CMD     : inout std_logic                     := '0';             --                       .hps_io_sdio_inst_CMD
		hps_io_hps_io_sdio_inst_D0      : inout std_logic                     := '0';             --                       .hps_io_sdio_inst_D0
		hps_io_hps_io_sdio_inst_D1      : inout std_logic                     := '0';             --                       .hps_io_sdio_inst_D1
		hps_io_hps_io_sdio_inst_CLK     : out   std_logic;                                        --                       .hps_io_sdio_inst_CLK
		hps_io_hps_io_sdio_inst_D2      : inout std_logic                     := '0';             --                       .hps_io_sdio_inst_D2
		hps_io_hps_io_sdio_inst_D3      : inout std_logic                     := '0';             --                       .hps_io_sdio_inst_D3
		hps_io_hps_io_usb1_inst_D0      : inout std_logic                     := '0';             --                       .hps_io_usb1_inst_D0
		hps_io_hps_io_usb1_inst_D1      : inout std_logic                     := '0';             --                       .hps_io_usb1_inst_D1
		hps_io_hps_io_usb1_inst_D2      : inout std_logic                     := '0';             --                       .hps_io_usb1_inst_D2
		hps_io_hps_io_usb1_inst_D3      : inout std_logic                     := '0';             --                       .hps_io_usb1_inst_D3
		hps_io_hps_io_usb1_inst_D4      : inout std_logic                     := '0';             --                       .hps_io_usb1_inst_D4
		hps_io_hps_io_usb1_inst_D5      : inout std_logic                     := '0';             --                       .hps_io_usb1_inst_D5
		hps_io_hps_io_usb1_inst_D6      : inout std_logic                     := '0';             --                       .hps_io_usb1_inst_D6
		hps_io_hps_io_usb1_inst_D7      : inout std_logic                     := '0';             --                       .hps_io_usb1_inst_D7
		hps_io_hps_io_usb1_inst_CLK     : in    std_logic                     := '0';             --                       .hps_io_usb1_inst_CLK
		hps_io_hps_io_usb1_inst_STP     : out   std_logic;                                        --                       .hps_io_usb1_inst_STP
		hps_io_hps_io_usb1_inst_DIR     : in    std_logic                     := '0';             --                       .hps_io_usb1_inst_DIR
		hps_io_hps_io_usb1_inst_NXT     : in    std_logic                     := '0';             --                       .hps_io_usb1_inst_NXT
		hps_io_hps_io_spim1_inst_CLK    : out   std_logic;                                        --                       .hps_io_spim1_inst_CLK
		hps_io_hps_io_spim1_inst_MOSI   : out   std_logic;                                        --                       .hps_io_spim1_inst_MOSI
		hps_io_hps_io_spim1_inst_MISO   : in    std_logic                     := '0';             --                       .hps_io_spim1_inst_MISO
		hps_io_hps_io_spim1_inst_SS0    : out   std_logic;                                        --                       .hps_io_spim1_inst_SS0
		hps_io_hps_io_uart0_inst_RX     : in    std_logic                     := '0';             --                       .hps_io_uart0_inst_RX
		hps_io_hps_io_uart0_inst_TX     : out   std_logic;                                        --                       .hps_io_uart0_inst_TX
		hps_io_hps_io_i2c1_inst_SDA     : inout std_logic                     := '0';             --                       .hps_io_i2c1_inst_SDA
		hps_io_hps_io_i2c1_inst_SCL     : inout std_logic                     := '0';             --                       .hps_io_i2c1_inst_SCL
		hps_io_hps_io_gpio_inst_GPIO09  : inout std_logic                     := '0';             --                       .hps_io_gpio_inst_GPIO09
		hps_io_hps_io_gpio_inst_GPIO35  : inout std_logic                     := '0';             --                       .hps_io_gpio_inst_GPIO35
		hps_io_hps_io_gpio_inst_GPIO40  : inout std_logic                     := '0';             --                       .hps_io_gpio_inst_GPIO40
		hps_io_hps_io_gpio_inst_GPIO53  : inout std_logic                     := '0';             --                       .hps_io_gpio_inst_GPIO53
		hps_io_hps_io_gpio_inst_GPIO54  : inout std_logic                     := '0';             --                       .hps_io_gpio_inst_GPIO54
		hps_io_hps_io_gpio_inst_GPIO61  : inout std_logic                     := '0';             --                       .hps_io_gpio_inst_GPIO61
		hps_spim0_txd                   : out   std_logic;                                        --              hps_spim0.txd
		hps_spim0_rxd                   : in    std_logic                     := '0';             --                       .rxd
		hps_spim0_ss_in_n               : in    std_logic                     := '0';             --                       .ss_in_n
		hps_spim0_ssi_oe_n              : out   std_logic;                                        --                       .ssi_oe_n
		hps_spim0_ss_0_n                : out   std_logic;                                        --                       .ss_0_n
		hps_spim0_ss_1_n                : out   std_logic;                                        --                       .ss_1_n
		hps_spim0_ss_2_n                : out   std_logic;                                        --                       .ss_2_n
		hps_spim0_ss_3_n                : out   std_logic;                                        --                       .ss_3_n
		hps_spim0_sclk_out_clk          : out   std_logic;                                        --     hps_spim0_sclk_out.clk
		memory_mem_a                    : out   std_logic_vector(14 downto 0);                    --                 memory.mem_a
		memory_mem_ba                   : out   std_logic_vector(2 downto 0);                     --                       .mem_ba
		memory_mem_ck                   : out   std_logic;                                        --                       .mem_ck
		memory_mem_ck_n                 : out   std_logic;                                        --                       .mem_ck_n
		memory_mem_cke                  : out   std_logic;                                        --                       .mem_cke
		memory_mem_cs_n                 : out   std_logic;                                        --                       .mem_cs_n
		memory_mem_ras_n                : out   std_logic;                                        --                       .mem_ras_n
		memory_mem_cas_n                : out   std_logic;                                        --                       .mem_cas_n
		memory_mem_we_n                 : out   std_logic;                                        --                       .mem_we_n
		memory_mem_reset_n              : out   std_logic;                                        --                       .mem_reset_n
		memory_mem_dq                   : inout std_logic_vector(31 downto 0) := (others => '0'); --                       .mem_dq
		memory_mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => '0'); --                       .mem_dqs
		memory_mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => '0'); --                       .mem_dqs_n
		memory_mem_odt                  : out   std_logic;                                        --                       .mem_odt
		memory_mem_dm                   : out   std_logic_vector(3 downto 0);                     --                       .mem_dm
		memory_oct_rzqin                : in    std_logic                     := '0'              --                       .oct_rzqin
	);
end entity soc_system_passthrough;

architecture rtl of soc_system_passthrough is
	component pitchshiftprocessor is
		port (
			reset                    : in  std_logic                     := 'X';             -- reset
			avalon_mm_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			avalon_mm_read           : in  std_logic                     := 'X';             -- read
			avalon_mm_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			avalon_mm_write          : in  std_logic                     := 'X';             -- write
			avalon_mm_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			clk                      : in  std_logic                     := 'X';             -- clk
			avalon_st_sink_channel   : in  std_logic                     := 'X';             -- channel
			avalon_st_sink_data      : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			avalon_st_sink_valid     : in  std_logic                     := 'X';             -- valid
			avalon_st_source_channel : out std_logic;                                        -- channel
			avalon_st_source_data    : out std_logic_vector(23 downto 0);                    -- data
			avalon_st_source_valid   : out std_logic                                         -- valid
		);
	end component pitchshiftprocessor;

	component soc_system_passthrough_ad1939_subsystem is
		port (
			ad1939_physical_asdata2     : in  std_logic                     := 'X';             -- asdata2
			ad1939_physical_dsdata1     : out std_logic;                                        -- dsdata1
			ad1939_physical_dbclk       : out std_logic;                                        -- dbclk
			ad1939_physical_dlrclk      : out std_logic;                                        -- dlrclk
			ad1939_physical_abclk_clk   : in  std_logic                     := 'X';             -- clk
			ad1939_physical_alrclk_clk  : in  std_logic                     := 'X';             -- clk
			ad1939_physical_mclk_clk    : in  std_logic                     := 'X';             -- clk
			audio_fabric_system_clk_clk : out std_logic;                                        -- clk
			from_line_in_data           : out std_logic_vector(23 downto 0);                    -- data
			from_line_in_channel        : out std_logic;                                        -- channel
			from_line_in_valid          : out std_logic;                                        -- valid
			subsystem_reset_reset       : in  std_logic                     := 'X';             -- reset
			to_headphone_out_data       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			to_headphone_out_channel    : in  std_logic                     := 'X';             -- channel
			to_headphone_out_valid      : in  std_logic                     := 'X'              -- valid
		);
	end component soc_system_passthrough_ad1939_subsystem;

	component soc_system_passthrough_audio_mini_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component soc_system_passthrough_audio_mini_leds;

	component soc_system_passthrough_clk_reset_inputs is
		port (
			fabric_reset_in_reset          : in  std_logic := 'X'; -- reset
			fabric_reset_out_reset         : out std_logic;        -- reset
			hps_and_fabric_reset_in_reset  : in  std_logic := 'X'; -- reset
			hps_and_fabric_reset_out_reset : out std_logic;        -- reset
			hps_clk_in_clk                 : in  std_logic := 'X'; -- clk
			hps_clk_out_clk                : out std_logic         -- clk
		);
	end component soc_system_passthrough_clk_reset_inputs;

	component soc_system_passthrough_de10_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component soc_system_passthrough_de10_leds;

	component soc_system_passthrough_hps is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			f2h_cold_rst_req_n       : in    std_logic                     := 'X';             -- reset_n
			spim0_txd                : out   std_logic;                                        -- txd
			spim0_rxd                : in    std_logic                     := 'X';             -- rxd
			spim0_ss_in_n            : in    std_logic                     := 'X';             -- ss_in_n
			spim0_ssi_oe_n           : out   std_logic;                                        -- ssi_oe_n
			spim0_ss_0_n             : out   std_logic;                                        -- ss_0_n
			spim0_ss_1_n             : out   std_logic;                                        -- ss_1_n
			spim0_ss_2_n             : out   std_logic;                                        -- ss_2_n
			spim0_ss_3_n             : out   std_logic;                                        -- ss_3_n
			spim0_sclk_out           : out   std_logic;                                        -- clk
			i2c0_scl                 : in    std_logic                     := 'X';             -- clk
			i2c0_out_clk             : out   std_logic;                                        -- clk
			i2c0_out_data            : out   std_logic;                                        -- out_data
			i2c0_sda                 : in    std_logic                     := 'X';             -- sda
			mem_a                    : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                   : out   std_logic;                                        -- mem_ck
			mem_ck_n                 : out   std_logic;                                        -- mem_ck_n
			mem_cke                  : out   std_logic;                                        -- mem_cke
			mem_cs_n                 : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                : out   std_logic;                                        -- mem_cas_n
			mem_we_n                 : out   std_logic;                                        -- mem_we_n
			mem_reset_n              : out   std_logic;                                        -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                        -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin                : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                        -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     : out   std_logic;                                        -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    : out   std_logic;                                        -- hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   : out   std_logic;                                        -- hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   : in    std_logic                     := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    : out   std_logic;                                        -- hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                        -- hps_io_uart0_inst_TX
			hps_io_i2c1_inst_SDA     : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO53  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO61
			h2f_rst_n                : out   std_logic;                                        -- reset_n
			h2f_lw_axi_clk           : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY           : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                        -- wlast
			h2f_lw_WVALID            : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY            : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                        -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY           : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic                                         -- rready
		);
	end component soc_system_passthrough_hps;

	component soc_system_passthrough_jtag_master is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component soc_system_passthrough_jtag_master;

	component soc_system_passthrough_system_id is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component soc_system_passthrough_system_id;

	component soc_system_passthrough_mm_interconnect_0 is
		port (
			hps_h2f_lw_axi_master_awid                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_h2f_lw_axi_master_awaddr                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_h2f_lw_axi_master_awlen                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_h2f_lw_axi_master_awsize                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_h2f_lw_axi_master_awburst                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_h2f_lw_axi_master_awlock                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_h2f_lw_axi_master_awcache                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_h2f_lw_axi_master_awprot                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_h2f_lw_axi_master_awvalid                     : in  std_logic                     := 'X';             -- awvalid
			hps_h2f_lw_axi_master_awready                     : out std_logic;                                        -- awready
			hps_h2f_lw_axi_master_wid                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_h2f_lw_axi_master_wdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_h2f_lw_axi_master_wstrb                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_h2f_lw_axi_master_wlast                       : in  std_logic                     := 'X';             -- wlast
			hps_h2f_lw_axi_master_wvalid                      : in  std_logic                     := 'X';             -- wvalid
			hps_h2f_lw_axi_master_wready                      : out std_logic;                                        -- wready
			hps_h2f_lw_axi_master_bid                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_h2f_lw_axi_master_bresp                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_h2f_lw_axi_master_bvalid                      : out std_logic;                                        -- bvalid
			hps_h2f_lw_axi_master_bready                      : in  std_logic                     := 'X';             -- bready
			hps_h2f_lw_axi_master_arid                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_h2f_lw_axi_master_araddr                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_h2f_lw_axi_master_arlen                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_h2f_lw_axi_master_arsize                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_h2f_lw_axi_master_arburst                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_h2f_lw_axi_master_arlock                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_h2f_lw_axi_master_arcache                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_h2f_lw_axi_master_arprot                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_h2f_lw_axi_master_arvalid                     : in  std_logic                     := 'X';             -- arvalid
			hps_h2f_lw_axi_master_arready                     : out std_logic;                                        -- arready
			hps_h2f_lw_axi_master_rid                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_h2f_lw_axi_master_rdata                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_h2f_lw_axi_master_rresp                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_h2f_lw_axi_master_rlast                       : out std_logic;                                        -- rlast
			hps_h2f_lw_axi_master_rvalid                      : out std_logic;                                        -- rvalid
			hps_h2f_lw_axi_master_rready                      : in  std_logic                     := 'X';             -- rready
			ad1939_subsystem_audio_fabric_system_clk_clk      : in  std_logic                     := 'X';             -- clk
			clk_reset_inputs_hps_clk_out_clk                  : in  std_logic                     := 'X';             -- clk
			audio_mini_leds_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			jtag_master_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			Pitch_Shift_0_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			system_id_reset_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			jtag_master_master_address                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			jtag_master_master_waitrequest                    : out std_logic;                                        -- waitrequest
			jtag_master_master_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_master_master_read                           : in  std_logic                     := 'X';             -- read
			jtag_master_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_master_master_readdatavalid                  : out std_logic;                                        -- readdatavalid
			jtag_master_master_write                          : in  std_logic                     := 'X';             -- write
			jtag_master_master_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			audio_mini_leds_s1_address                        : out std_logic_vector(1 downto 0);                     -- address
			audio_mini_leds_s1_write                          : out std_logic;                                        -- write
			audio_mini_leds_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_mini_leds_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			audio_mini_leds_s1_chipselect                     : out std_logic;                                        -- chipselect
			de10_leds_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			de10_leds_s1_write                                : out std_logic;                                        -- write
			de10_leds_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			de10_leds_s1_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			de10_leds_s1_chipselect                           : out std_logic;                                        -- chipselect
			Pitch_Shift_0_avalon_mm_address                   : out std_logic_vector(1 downto 0);                     -- address
			Pitch_Shift_0_avalon_mm_write                     : out std_logic;                                        -- write
			Pitch_Shift_0_avalon_mm_read                      : out std_logic;                                        -- read
			Pitch_Shift_0_avalon_mm_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Pitch_Shift_0_avalon_mm_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			system_id_control_slave_address                   : out std_logic_vector(0 downto 0);                     -- address
			system_id_control_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component soc_system_passthrough_mm_interconnect_0;

	component soc_system_passthrough_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_passthrough_rst_controller;

	component soc_system_passthrough_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_passthrough_rst_controller_002;

	signal pitch_shift_0_avalon_streaming_source_valid               : std_logic;                     -- Pitch_Shift_0:avalon_st_source_valid -> ad1939_subsystem:to_headphone_out_valid
	signal pitch_shift_0_avalon_streaming_source_data                : std_logic_vector(23 downto 0); -- Pitch_Shift_0:avalon_st_source_data -> ad1939_subsystem:to_headphone_out_data
	signal pitch_shift_0_avalon_streaming_source_channel             : std_logic;                     -- Pitch_Shift_0:avalon_st_source_channel -> ad1939_subsystem:to_headphone_out_channel
	signal ad1939_subsystem_from_line_in_valid                       : std_logic;                     -- ad1939_subsystem:from_line_in_valid -> Pitch_Shift_0:avalon_st_sink_valid
	signal ad1939_subsystem_from_line_in_data                        : std_logic_vector(23 downto 0); -- ad1939_subsystem:from_line_in_data -> Pitch_Shift_0:avalon_st_sink_data
	signal ad1939_subsystem_from_line_in_channel                     : std_logic;                     -- ad1939_subsystem:from_line_in_channel -> Pitch_Shift_0:avalon_st_sink_channel
	signal ad1939_subsystem_audio_fabric_system_clk_clk              : std_logic;                     -- ad1939_subsystem:audio_fabric_system_clk_clk -> [Pitch_Shift_0:clk, mm_interconnect_0:ad1939_subsystem_audio_fabric_system_clk_clk, rst_controller:clk]
	signal clk_reset_inputs_hps_clk_out_clk                          : std_logic;                     -- clk_reset_inputs:hps_clk_out_clk -> [audio_mini_leds:clk, de10_leds:clk, hps:h2f_lw_axi_clk, jtag_master:clk_clk, mm_interconnect_0:clk_reset_inputs_hps_clk_out_clk, rst_controller_002:clk, rst_controller_003:clk, system_id:clock]
	signal hps_h2f_reset_reset                                       : std_logic;                     -- hps:h2f_rst_n -> hps_h2f_reset_reset:in
	signal clk_reset_inputs_hps_and_fabric_reset_out_reset           : std_logic;                     -- clk_reset_inputs:hps_and_fabric_reset_out_reset -> [clk_reset_inputs_hps_and_fabric_reset_out_reset:in, rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	signal hps_h2f_lw_axi_master_awburst                             : std_logic_vector(1 downto 0);  -- hps:h2f_lw_AWBURST -> mm_interconnect_0:hps_h2f_lw_axi_master_awburst
	signal hps_h2f_lw_axi_master_arlen                               : std_logic_vector(3 downto 0);  -- hps:h2f_lw_ARLEN -> mm_interconnect_0:hps_h2f_lw_axi_master_arlen
	signal hps_h2f_lw_axi_master_wstrb                               : std_logic_vector(3 downto 0);  -- hps:h2f_lw_WSTRB -> mm_interconnect_0:hps_h2f_lw_axi_master_wstrb
	signal hps_h2f_lw_axi_master_wready                              : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_wready -> hps:h2f_lw_WREADY
	signal hps_h2f_lw_axi_master_rid                                 : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_h2f_lw_axi_master_rid -> hps:h2f_lw_RID
	signal hps_h2f_lw_axi_master_rready                              : std_logic;                     -- hps:h2f_lw_RREADY -> mm_interconnect_0:hps_h2f_lw_axi_master_rready
	signal hps_h2f_lw_axi_master_awlen                               : std_logic_vector(3 downto 0);  -- hps:h2f_lw_AWLEN -> mm_interconnect_0:hps_h2f_lw_axi_master_awlen
	signal hps_h2f_lw_axi_master_wid                                 : std_logic_vector(11 downto 0); -- hps:h2f_lw_WID -> mm_interconnect_0:hps_h2f_lw_axi_master_wid
	signal hps_h2f_lw_axi_master_arcache                             : std_logic_vector(3 downto 0);  -- hps:h2f_lw_ARCACHE -> mm_interconnect_0:hps_h2f_lw_axi_master_arcache
	signal hps_h2f_lw_axi_master_wvalid                              : std_logic;                     -- hps:h2f_lw_WVALID -> mm_interconnect_0:hps_h2f_lw_axi_master_wvalid
	signal hps_h2f_lw_axi_master_araddr                              : std_logic_vector(20 downto 0); -- hps:h2f_lw_ARADDR -> mm_interconnect_0:hps_h2f_lw_axi_master_araddr
	signal hps_h2f_lw_axi_master_arprot                              : std_logic_vector(2 downto 0);  -- hps:h2f_lw_ARPROT -> mm_interconnect_0:hps_h2f_lw_axi_master_arprot
	signal hps_h2f_lw_axi_master_awprot                              : std_logic_vector(2 downto 0);  -- hps:h2f_lw_AWPROT -> mm_interconnect_0:hps_h2f_lw_axi_master_awprot
	signal hps_h2f_lw_axi_master_wdata                               : std_logic_vector(31 downto 0); -- hps:h2f_lw_WDATA -> mm_interconnect_0:hps_h2f_lw_axi_master_wdata
	signal hps_h2f_lw_axi_master_arvalid                             : std_logic;                     -- hps:h2f_lw_ARVALID -> mm_interconnect_0:hps_h2f_lw_axi_master_arvalid
	signal hps_h2f_lw_axi_master_awcache                             : std_logic_vector(3 downto 0);  -- hps:h2f_lw_AWCACHE -> mm_interconnect_0:hps_h2f_lw_axi_master_awcache
	signal hps_h2f_lw_axi_master_arid                                : std_logic_vector(11 downto 0); -- hps:h2f_lw_ARID -> mm_interconnect_0:hps_h2f_lw_axi_master_arid
	signal hps_h2f_lw_axi_master_arlock                              : std_logic_vector(1 downto 0);  -- hps:h2f_lw_ARLOCK -> mm_interconnect_0:hps_h2f_lw_axi_master_arlock
	signal hps_h2f_lw_axi_master_awlock                              : std_logic_vector(1 downto 0);  -- hps:h2f_lw_AWLOCK -> mm_interconnect_0:hps_h2f_lw_axi_master_awlock
	signal hps_h2f_lw_axi_master_awaddr                              : std_logic_vector(20 downto 0); -- hps:h2f_lw_AWADDR -> mm_interconnect_0:hps_h2f_lw_axi_master_awaddr
	signal hps_h2f_lw_axi_master_bresp                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_h2f_lw_axi_master_bresp -> hps:h2f_lw_BRESP
	signal hps_h2f_lw_axi_master_arready                             : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_arready -> hps:h2f_lw_ARREADY
	signal hps_h2f_lw_axi_master_rdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:hps_h2f_lw_axi_master_rdata -> hps:h2f_lw_RDATA
	signal hps_h2f_lw_axi_master_awready                             : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_awready -> hps:h2f_lw_AWREADY
	signal hps_h2f_lw_axi_master_arburst                             : std_logic_vector(1 downto 0);  -- hps:h2f_lw_ARBURST -> mm_interconnect_0:hps_h2f_lw_axi_master_arburst
	signal hps_h2f_lw_axi_master_arsize                              : std_logic_vector(2 downto 0);  -- hps:h2f_lw_ARSIZE -> mm_interconnect_0:hps_h2f_lw_axi_master_arsize
	signal hps_h2f_lw_axi_master_bready                              : std_logic;                     -- hps:h2f_lw_BREADY -> mm_interconnect_0:hps_h2f_lw_axi_master_bready
	signal hps_h2f_lw_axi_master_rlast                               : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_rlast -> hps:h2f_lw_RLAST
	signal hps_h2f_lw_axi_master_wlast                               : std_logic;                     -- hps:h2f_lw_WLAST -> mm_interconnect_0:hps_h2f_lw_axi_master_wlast
	signal hps_h2f_lw_axi_master_rresp                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_h2f_lw_axi_master_rresp -> hps:h2f_lw_RRESP
	signal hps_h2f_lw_axi_master_awid                                : std_logic_vector(11 downto 0); -- hps:h2f_lw_AWID -> mm_interconnect_0:hps_h2f_lw_axi_master_awid
	signal hps_h2f_lw_axi_master_bid                                 : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_h2f_lw_axi_master_bid -> hps:h2f_lw_BID
	signal hps_h2f_lw_axi_master_bvalid                              : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_bvalid -> hps:h2f_lw_BVALID
	signal hps_h2f_lw_axi_master_awsize                              : std_logic_vector(2 downto 0);  -- hps:h2f_lw_AWSIZE -> mm_interconnect_0:hps_h2f_lw_axi_master_awsize
	signal hps_h2f_lw_axi_master_awvalid                             : std_logic;                     -- hps:h2f_lw_AWVALID -> mm_interconnect_0:hps_h2f_lw_axi_master_awvalid
	signal hps_h2f_lw_axi_master_rvalid                              : std_logic;                     -- mm_interconnect_0:hps_h2f_lw_axi_master_rvalid -> hps:h2f_lw_RVALID
	signal jtag_master_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_master_master_readdata -> jtag_master:master_readdata
	signal jtag_master_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:jtag_master_master_waitrequest -> jtag_master:master_waitrequest
	signal jtag_master_master_address                                : std_logic_vector(31 downto 0); -- jtag_master:master_address -> mm_interconnect_0:jtag_master_master_address
	signal jtag_master_master_read                                   : std_logic;                     -- jtag_master:master_read -> mm_interconnect_0:jtag_master_master_read
	signal jtag_master_master_byteenable                             : std_logic_vector(3 downto 0);  -- jtag_master:master_byteenable -> mm_interconnect_0:jtag_master_master_byteenable
	signal jtag_master_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:jtag_master_master_readdatavalid -> jtag_master:master_readdatavalid
	signal jtag_master_master_write                                  : std_logic;                     -- jtag_master:master_write -> mm_interconnect_0:jtag_master_master_write
	signal jtag_master_master_writedata                              : std_logic_vector(31 downto 0); -- jtag_master:master_writedata -> mm_interconnect_0:jtag_master_master_writedata
	signal mm_interconnect_0_pitch_shift_0_avalon_mm_readdata        : std_logic_vector(31 downto 0); -- Pitch_Shift_0:avalon_mm_readdata -> mm_interconnect_0:Pitch_Shift_0_avalon_mm_readdata
	signal mm_interconnect_0_pitch_shift_0_avalon_mm_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Pitch_Shift_0_avalon_mm_address -> Pitch_Shift_0:avalon_mm_address
	signal mm_interconnect_0_pitch_shift_0_avalon_mm_read            : std_logic;                     -- mm_interconnect_0:Pitch_Shift_0_avalon_mm_read -> Pitch_Shift_0:avalon_mm_read
	signal mm_interconnect_0_pitch_shift_0_avalon_mm_write           : std_logic;                     -- mm_interconnect_0:Pitch_Shift_0_avalon_mm_write -> Pitch_Shift_0:avalon_mm_write
	signal mm_interconnect_0_pitch_shift_0_avalon_mm_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:Pitch_Shift_0_avalon_mm_writedata -> Pitch_Shift_0:avalon_mm_writedata
	signal mm_interconnect_0_system_id_control_slave_readdata        : std_logic_vector(31 downto 0); -- system_id:readdata -> mm_interconnect_0:system_id_control_slave_readdata
	signal mm_interconnect_0_system_id_control_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:system_id_control_slave_address -> system_id:address
	signal mm_interconnect_0_audio_mini_leds_s1_chipselect           : std_logic;                     -- mm_interconnect_0:audio_mini_leds_s1_chipselect -> audio_mini_leds:chipselect
	signal mm_interconnect_0_audio_mini_leds_s1_readdata             : std_logic_vector(31 downto 0); -- audio_mini_leds:readdata -> mm_interconnect_0:audio_mini_leds_s1_readdata
	signal mm_interconnect_0_audio_mini_leds_s1_address              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_mini_leds_s1_address -> audio_mini_leds:address
	signal mm_interconnect_0_audio_mini_leds_s1_write                : std_logic;                     -- mm_interconnect_0:audio_mini_leds_s1_write -> mm_interconnect_0_audio_mini_leds_s1_write:in
	signal mm_interconnect_0_audio_mini_leds_s1_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_mini_leds_s1_writedata -> audio_mini_leds:writedata
	signal mm_interconnect_0_de10_leds_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:de10_leds_s1_chipselect -> de10_leds:chipselect
	signal mm_interconnect_0_de10_leds_s1_readdata                   : std_logic_vector(31 downto 0); -- de10_leds:readdata -> mm_interconnect_0:de10_leds_s1_readdata
	signal mm_interconnect_0_de10_leds_s1_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:de10_leds_s1_address -> de10_leds:address
	signal mm_interconnect_0_de10_leds_s1_write                      : std_logic;                     -- mm_interconnect_0:de10_leds_s1_write -> mm_interconnect_0_de10_leds_s1_write:in
	signal mm_interconnect_0_de10_leds_s1_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:de10_leds_s1_writedata -> de10_leds:writedata
	signal rst_controller_reset_out_reset                            : std_logic;                     -- rst_controller:reset_out -> [Pitch_Shift_0:reset, mm_interconnect_0:Pitch_Shift_0_reset_reset_bridge_in_reset_reset]
	signal clk_reset_inputs_fabric_reset_out_reset                   : std_logic;                     -- clk_reset_inputs:fabric_reset_out_reset -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal rst_controller_001_reset_out_reset                        : std_logic;                     -- rst_controller_001:reset_out -> ad1939_subsystem:subsystem_reset_reset
	signal rst_controller_002_reset_out_reset                        : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:audio_mini_leds_reset_reset_bridge_in_reset_reset, rst_controller_002_reset_out_reset:in]
	signal rst_controller_003_reset_out_reset                        : std_logic;                     -- rst_controller_003:reset_out -> [mm_interconnect_0:jtag_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:system_id_reset_reset_bridge_in_reset_reset, rst_controller_003_reset_out_reset:in]
	signal hps_h2f_reset_reset_ports_inv                             : std_logic;                     -- hps_h2f_reset_reset:inv -> [jtag_master:clk_reset_reset, rst_controller_003:reset_in0]
	signal clk_reset_inputs_hps_and_fabric_reset_out_reset_ports_inv : std_logic;                     -- clk_reset_inputs_hps_and_fabric_reset_out_reset:inv -> hps:f2h_cold_rst_req_n
	signal mm_interconnect_0_audio_mini_leds_s1_write_ports_inv      : std_logic;                     -- mm_interconnect_0_audio_mini_leds_s1_write:inv -> audio_mini_leds:write_n
	signal mm_interconnect_0_de10_leds_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_0_de10_leds_s1_write:inv -> de10_leds:write_n
	signal rst_controller_002_reset_out_reset_ports_inv              : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> [audio_mini_leds:reset_n, de10_leds:reset_n]
	signal rst_controller_003_reset_out_reset_ports_inv              : std_logic;                     -- rst_controller_003_reset_out_reset:inv -> system_id:reset_n

begin

	pitch_shift_0 : component pitchshiftprocessor
		port map (
			reset                    => rst_controller_reset_out_reset,                      --                   reset.reset
			avalon_mm_address        => mm_interconnect_0_pitch_shift_0_avalon_mm_address,   --               avalon_mm.address
			avalon_mm_read           => mm_interconnect_0_pitch_shift_0_avalon_mm_read,      --                        .read
			avalon_mm_readdata       => mm_interconnect_0_pitch_shift_0_avalon_mm_readdata,  --                        .readdata
			avalon_mm_write          => mm_interconnect_0_pitch_shift_0_avalon_mm_write,     --                        .write
			avalon_mm_writedata      => mm_interconnect_0_pitch_shift_0_avalon_mm_writedata, --                        .writedata
			clk                      => ad1939_subsystem_audio_fabric_system_clk_clk,        --                   clock.clk
			avalon_st_sink_channel   => ad1939_subsystem_from_line_in_channel,               --   avalon_streaming_sink.channel
			avalon_st_sink_data      => ad1939_subsystem_from_line_in_data,                  --                        .data
			avalon_st_sink_valid     => ad1939_subsystem_from_line_in_valid,                 --                        .valid
			avalon_st_source_channel => pitch_shift_0_avalon_streaming_source_channel,       -- avalon_streaming_source.channel
			avalon_st_source_data    => pitch_shift_0_avalon_streaming_source_data,          --                        .data
			avalon_st_source_valid   => pitch_shift_0_avalon_streaming_source_valid          --                        .valid
		);

	ad1939_subsystem : component soc_system_passthrough_ad1939_subsystem
		port map (
			ad1939_physical_asdata2     => ad1939_physical_asdata2,                       --         ad1939_physical.asdata2
			ad1939_physical_dsdata1     => ad1939_physical_dsdata1,                       --                        .dsdata1
			ad1939_physical_dbclk       => ad1939_physical_dbclk,                         --                        .dbclk
			ad1939_physical_dlrclk      => ad1939_physical_dlrclk,                        --                        .dlrclk
			ad1939_physical_abclk_clk   => ad1939_physical_abclk_clk,                     --   ad1939_physical_abclk.clk
			ad1939_physical_alrclk_clk  => ad1939_physical_alrclk_clk,                    --  ad1939_physical_alrclk.clk
			ad1939_physical_mclk_clk    => ad1939_physical_mclk_clk,                      --    ad1939_physical_mclk.clk
			audio_fabric_system_clk_clk => ad1939_subsystem_audio_fabric_system_clk_clk,  -- audio_fabric_system_clk.clk
			from_line_in_data           => ad1939_subsystem_from_line_in_data,            --            from_line_in.data
			from_line_in_channel        => ad1939_subsystem_from_line_in_channel,         --                        .channel
			from_line_in_valid          => ad1939_subsystem_from_line_in_valid,           --                        .valid
			subsystem_reset_reset       => rst_controller_001_reset_out_reset,            --         subsystem_reset.reset
			to_headphone_out_data       => pitch_shift_0_avalon_streaming_source_data,    --        to_headphone_out.data
			to_headphone_out_channel    => pitch_shift_0_avalon_streaming_source_channel, --                        .channel
			to_headphone_out_valid      => pitch_shift_0_avalon_streaming_source_valid    --                        .valid
		);

	audio_mini_leds : component soc_system_passthrough_audio_mini_leds
		port map (
			clk        => clk_reset_inputs_hps_clk_out_clk,                     --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_audio_mini_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_audio_mini_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_audio_mini_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_audio_mini_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_audio_mini_leds_s1_readdata,        --                    .readdata
			out_port   => audio_mini_leds_export                                -- external_connection.export
		);

	clk_reset_inputs : component soc_system_passthrough_clk_reset_inputs
		port map (
			fabric_reset_in_reset          => fabric_reset_reset,                              --          fabric_reset_in.reset
			fabric_reset_out_reset         => clk_reset_inputs_fabric_reset_out_reset,         --         fabric_reset_out.reset
			hps_and_fabric_reset_in_reset  => hps_and_fabric_reset_reset,                      --  hps_and_fabric_reset_in.reset
			hps_and_fabric_reset_out_reset => clk_reset_inputs_hps_and_fabric_reset_out_reset, -- hps_and_fabric_reset_out.reset
			hps_clk_in_clk                 => hps_clk_clk,                                     --               hps_clk_in.clk
			hps_clk_out_clk                => clk_reset_inputs_hps_clk_out_clk                 --              hps_clk_out.clk
		);

	de10_leds : component soc_system_passthrough_de10_leds
		port map (
			clk        => clk_reset_inputs_hps_clk_out_clk,               --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_de10_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_de10_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_de10_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_de10_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_de10_leds_s1_readdata,        --                    .readdata
			out_port   => de10_leds_export                                -- external_connection.export
		);

	hps : component soc_system_passthrough_hps
		generic map (
			F2S_Width => 0,
			S2F_Width => 0
		)
		port map (
			f2h_cold_rst_req_n       => clk_reset_inputs_hps_and_fabric_reset_out_reset_ports_inv, -- f2h_cold_reset_req.reset_n
			spim0_txd                => hps_spim0_txd,                                             --              spim0.txd
			spim0_rxd                => hps_spim0_rxd,                                             --                   .rxd
			spim0_ss_in_n            => hps_spim0_ss_in_n,                                         --                   .ss_in_n
			spim0_ssi_oe_n           => hps_spim0_ssi_oe_n,                                        --                   .ssi_oe_n
			spim0_ss_0_n             => hps_spim0_ss_0_n,                                          --                   .ss_0_n
			spim0_ss_1_n             => hps_spim0_ss_1_n,                                          --                   .ss_1_n
			spim0_ss_2_n             => hps_spim0_ss_2_n,                                          --                   .ss_2_n
			spim0_ss_3_n             => hps_spim0_ss_3_n,                                          --                   .ss_3_n
			spim0_sclk_out           => hps_spim0_sclk_out_clk,                                    --     spim0_sclk_out.clk
			i2c0_scl                 => hps_i2c0_scl_in_clk,                                       --        i2c0_scl_in.clk
			i2c0_out_clk             => hps_i2c0_clk_clk,                                          --           i2c0_clk.clk
			i2c0_out_data            => hps_i2c0_out_data,                                         --               i2c0.out_data
			i2c0_sda                 => hps_i2c0_sda,                                              --                   .sda
			mem_a                    => memory_mem_a,                                              --             memory.mem_a
			mem_ba                   => memory_mem_ba,                                             --                   .mem_ba
			mem_ck                   => memory_mem_ck,                                             --                   .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                                           --                   .mem_ck_n
			mem_cke                  => memory_mem_cke,                                            --                   .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                                           --                   .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                                          --                   .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                                          --                   .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                                           --                   .mem_we_n
			mem_reset_n              => memory_mem_reset_n,                                        --                   .mem_reset_n
			mem_dq                   => memory_mem_dq,                                             --                   .mem_dq
			mem_dqs                  => memory_mem_dqs,                                            --                   .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                                          --                   .mem_dqs_n
			mem_odt                  => memory_mem_odt,                                            --                   .mem_odt
			mem_dm                   => memory_mem_dm,                                             --                   .mem_dm
			oct_rzqin                => memory_oct_rzqin,                                          --                   .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_io_hps_io_emac1_inst_TX_CLK,                           --             hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_io_hps_io_emac1_inst_TXD0,                             --                   .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_io_hps_io_emac1_inst_TXD1,                             --                   .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_io_hps_io_emac1_inst_TXD2,                             --                   .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_io_hps_io_emac1_inst_TXD3,                             --                   .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_io_hps_io_emac1_inst_RXD0,                             --                   .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_io_hps_io_emac1_inst_MDIO,                             --                   .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_io_hps_io_emac1_inst_MDC,                              --                   .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_io_hps_io_emac1_inst_RX_CTL,                           --                   .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_io_hps_io_emac1_inst_TX_CTL,                           --                   .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_io_hps_io_emac1_inst_RX_CLK,                           --                   .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_io_hps_io_emac1_inst_RXD1,                             --                   .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_io_hps_io_emac1_inst_RXD2,                             --                   .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_io_hps_io_emac1_inst_RXD3,                             --                   .hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     => hps_io_hps_io_sdio_inst_CMD,                               --                   .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_io_hps_io_sdio_inst_D0,                                --                   .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_io_hps_io_sdio_inst_D1,                                --                   .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_io_hps_io_sdio_inst_CLK,                               --                   .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_io_hps_io_sdio_inst_D2,                                --                   .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_io_hps_io_sdio_inst_D3,                                --                   .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      => hps_io_hps_io_usb1_inst_D0,                                --                   .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      => hps_io_hps_io_usb1_inst_D1,                                --                   .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      => hps_io_hps_io_usb1_inst_D2,                                --                   .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      => hps_io_hps_io_usb1_inst_D3,                                --                   .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      => hps_io_hps_io_usb1_inst_D4,                                --                   .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      => hps_io_hps_io_usb1_inst_D5,                                --                   .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      => hps_io_hps_io_usb1_inst_D6,                                --                   .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      => hps_io_hps_io_usb1_inst_D7,                                --                   .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     => hps_io_hps_io_usb1_inst_CLK,                               --                   .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     => hps_io_hps_io_usb1_inst_STP,                               --                   .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     => hps_io_hps_io_usb1_inst_DIR,                               --                   .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     => hps_io_hps_io_usb1_inst_NXT,                               --                   .hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    => hps_io_hps_io_spim1_inst_CLK,                              --                   .hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   => hps_io_hps_io_spim1_inst_MOSI,                             --                   .hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   => hps_io_hps_io_spim1_inst_MISO,                             --                   .hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    => hps_io_hps_io_spim1_inst_SS0,                              --                   .hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     => hps_io_hps_io_uart0_inst_RX,                               --                   .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_io_hps_io_uart0_inst_TX,                               --                   .hps_io_uart0_inst_TX
			hps_io_i2c1_inst_SDA     => hps_io_hps_io_i2c1_inst_SDA,                               --                   .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     => hps_io_hps_io_i2c1_inst_SCL,                               --                   .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  => hps_io_hps_io_gpio_inst_GPIO09,                            --                   .hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  => hps_io_hps_io_gpio_inst_GPIO35,                            --                   .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  => hps_io_hps_io_gpio_inst_GPIO40,                            --                   .hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO53  => hps_io_hps_io_gpio_inst_GPIO53,                            --                   .hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  => hps_io_hps_io_gpio_inst_GPIO54,                            --                   .hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  => hps_io_hps_io_gpio_inst_GPIO61,                            --                   .hps_io_gpio_inst_GPIO61
			h2f_rst_n                => hps_h2f_reset_reset,                                       --          h2f_reset.reset_n
			h2f_lw_axi_clk           => clk_reset_inputs_hps_clk_out_clk,                          --   h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_h2f_lw_axi_master_awid,                                --  h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_h2f_lw_axi_master_awaddr,                              --                   .awaddr
			h2f_lw_AWLEN             => hps_h2f_lw_axi_master_awlen,                               --                   .awlen
			h2f_lw_AWSIZE            => hps_h2f_lw_axi_master_awsize,                              --                   .awsize
			h2f_lw_AWBURST           => hps_h2f_lw_axi_master_awburst,                             --                   .awburst
			h2f_lw_AWLOCK            => hps_h2f_lw_axi_master_awlock,                              --                   .awlock
			h2f_lw_AWCACHE           => hps_h2f_lw_axi_master_awcache,                             --                   .awcache
			h2f_lw_AWPROT            => hps_h2f_lw_axi_master_awprot,                              --                   .awprot
			h2f_lw_AWVALID           => hps_h2f_lw_axi_master_awvalid,                             --                   .awvalid
			h2f_lw_AWREADY           => hps_h2f_lw_axi_master_awready,                             --                   .awready
			h2f_lw_WID               => hps_h2f_lw_axi_master_wid,                                 --                   .wid
			h2f_lw_WDATA             => hps_h2f_lw_axi_master_wdata,                               --                   .wdata
			h2f_lw_WSTRB             => hps_h2f_lw_axi_master_wstrb,                               --                   .wstrb
			h2f_lw_WLAST             => hps_h2f_lw_axi_master_wlast,                               --                   .wlast
			h2f_lw_WVALID            => hps_h2f_lw_axi_master_wvalid,                              --                   .wvalid
			h2f_lw_WREADY            => hps_h2f_lw_axi_master_wready,                              --                   .wready
			h2f_lw_BID               => hps_h2f_lw_axi_master_bid,                                 --                   .bid
			h2f_lw_BRESP             => hps_h2f_lw_axi_master_bresp,                               --                   .bresp
			h2f_lw_BVALID            => hps_h2f_lw_axi_master_bvalid,                              --                   .bvalid
			h2f_lw_BREADY            => hps_h2f_lw_axi_master_bready,                              --                   .bready
			h2f_lw_ARID              => hps_h2f_lw_axi_master_arid,                                --                   .arid
			h2f_lw_ARADDR            => hps_h2f_lw_axi_master_araddr,                              --                   .araddr
			h2f_lw_ARLEN             => hps_h2f_lw_axi_master_arlen,                               --                   .arlen
			h2f_lw_ARSIZE            => hps_h2f_lw_axi_master_arsize,                              --                   .arsize
			h2f_lw_ARBURST           => hps_h2f_lw_axi_master_arburst,                             --                   .arburst
			h2f_lw_ARLOCK            => hps_h2f_lw_axi_master_arlock,                              --                   .arlock
			h2f_lw_ARCACHE           => hps_h2f_lw_axi_master_arcache,                             --                   .arcache
			h2f_lw_ARPROT            => hps_h2f_lw_axi_master_arprot,                              --                   .arprot
			h2f_lw_ARVALID           => hps_h2f_lw_axi_master_arvalid,                             --                   .arvalid
			h2f_lw_ARREADY           => hps_h2f_lw_axi_master_arready,                             --                   .arready
			h2f_lw_RID               => hps_h2f_lw_axi_master_rid,                                 --                   .rid
			h2f_lw_RDATA             => hps_h2f_lw_axi_master_rdata,                               --                   .rdata
			h2f_lw_RRESP             => hps_h2f_lw_axi_master_rresp,                               --                   .rresp
			h2f_lw_RLAST             => hps_h2f_lw_axi_master_rlast,                               --                   .rlast
			h2f_lw_RVALID            => hps_h2f_lw_axi_master_rvalid,                              --                   .rvalid
			h2f_lw_RREADY            => hps_h2f_lw_axi_master_rready                               --                   .rready
		);

	jtag_master : component soc_system_passthrough_jtag_master
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => clk_reset_inputs_hps_clk_out_clk, --          clk.clk
			clk_reset_reset      => hps_h2f_reset_reset_ports_inv,    --    clk_reset.reset
			master_address       => jtag_master_master_address,       --       master.address
			master_readdata      => jtag_master_master_readdata,      --             .readdata
			master_read          => jtag_master_master_read,          --             .read
			master_write         => jtag_master_master_write,         --             .write
			master_writedata     => jtag_master_master_writedata,     --             .writedata
			master_waitrequest   => jtag_master_master_waitrequest,   --             .waitrequest
			master_readdatavalid => jtag_master_master_readdatavalid, --             .readdatavalid
			master_byteenable    => jtag_master_master_byteenable,    --             .byteenable
			master_reset_reset   => open                              -- master_reset.reset
		);

	system_id : component soc_system_passthrough_system_id
		port map (
			clock    => clk_reset_inputs_hps_clk_out_clk,                     --           clk.clk
			reset_n  => rst_controller_003_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_system_id_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_system_id_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component soc_system_passthrough_mm_interconnect_0
		port map (
			hps_h2f_lw_axi_master_awid                        => hps_h2f_lw_axi_master_awid,                          --                       hps_h2f_lw_axi_master.awid
			hps_h2f_lw_axi_master_awaddr                      => hps_h2f_lw_axi_master_awaddr,                        --                                            .awaddr
			hps_h2f_lw_axi_master_awlen                       => hps_h2f_lw_axi_master_awlen,                         --                                            .awlen
			hps_h2f_lw_axi_master_awsize                      => hps_h2f_lw_axi_master_awsize,                        --                                            .awsize
			hps_h2f_lw_axi_master_awburst                     => hps_h2f_lw_axi_master_awburst,                       --                                            .awburst
			hps_h2f_lw_axi_master_awlock                      => hps_h2f_lw_axi_master_awlock,                        --                                            .awlock
			hps_h2f_lw_axi_master_awcache                     => hps_h2f_lw_axi_master_awcache,                       --                                            .awcache
			hps_h2f_lw_axi_master_awprot                      => hps_h2f_lw_axi_master_awprot,                        --                                            .awprot
			hps_h2f_lw_axi_master_awvalid                     => hps_h2f_lw_axi_master_awvalid,                       --                                            .awvalid
			hps_h2f_lw_axi_master_awready                     => hps_h2f_lw_axi_master_awready,                       --                                            .awready
			hps_h2f_lw_axi_master_wid                         => hps_h2f_lw_axi_master_wid,                           --                                            .wid
			hps_h2f_lw_axi_master_wdata                       => hps_h2f_lw_axi_master_wdata,                         --                                            .wdata
			hps_h2f_lw_axi_master_wstrb                       => hps_h2f_lw_axi_master_wstrb,                         --                                            .wstrb
			hps_h2f_lw_axi_master_wlast                       => hps_h2f_lw_axi_master_wlast,                         --                                            .wlast
			hps_h2f_lw_axi_master_wvalid                      => hps_h2f_lw_axi_master_wvalid,                        --                                            .wvalid
			hps_h2f_lw_axi_master_wready                      => hps_h2f_lw_axi_master_wready,                        --                                            .wready
			hps_h2f_lw_axi_master_bid                         => hps_h2f_lw_axi_master_bid,                           --                                            .bid
			hps_h2f_lw_axi_master_bresp                       => hps_h2f_lw_axi_master_bresp,                         --                                            .bresp
			hps_h2f_lw_axi_master_bvalid                      => hps_h2f_lw_axi_master_bvalid,                        --                                            .bvalid
			hps_h2f_lw_axi_master_bready                      => hps_h2f_lw_axi_master_bready,                        --                                            .bready
			hps_h2f_lw_axi_master_arid                        => hps_h2f_lw_axi_master_arid,                          --                                            .arid
			hps_h2f_lw_axi_master_araddr                      => hps_h2f_lw_axi_master_araddr,                        --                                            .araddr
			hps_h2f_lw_axi_master_arlen                       => hps_h2f_lw_axi_master_arlen,                         --                                            .arlen
			hps_h2f_lw_axi_master_arsize                      => hps_h2f_lw_axi_master_arsize,                        --                                            .arsize
			hps_h2f_lw_axi_master_arburst                     => hps_h2f_lw_axi_master_arburst,                       --                                            .arburst
			hps_h2f_lw_axi_master_arlock                      => hps_h2f_lw_axi_master_arlock,                        --                                            .arlock
			hps_h2f_lw_axi_master_arcache                     => hps_h2f_lw_axi_master_arcache,                       --                                            .arcache
			hps_h2f_lw_axi_master_arprot                      => hps_h2f_lw_axi_master_arprot,                        --                                            .arprot
			hps_h2f_lw_axi_master_arvalid                     => hps_h2f_lw_axi_master_arvalid,                       --                                            .arvalid
			hps_h2f_lw_axi_master_arready                     => hps_h2f_lw_axi_master_arready,                       --                                            .arready
			hps_h2f_lw_axi_master_rid                         => hps_h2f_lw_axi_master_rid,                           --                                            .rid
			hps_h2f_lw_axi_master_rdata                       => hps_h2f_lw_axi_master_rdata,                         --                                            .rdata
			hps_h2f_lw_axi_master_rresp                       => hps_h2f_lw_axi_master_rresp,                         --                                            .rresp
			hps_h2f_lw_axi_master_rlast                       => hps_h2f_lw_axi_master_rlast,                         --                                            .rlast
			hps_h2f_lw_axi_master_rvalid                      => hps_h2f_lw_axi_master_rvalid,                        --                                            .rvalid
			hps_h2f_lw_axi_master_rready                      => hps_h2f_lw_axi_master_rready,                        --                                            .rready
			ad1939_subsystem_audio_fabric_system_clk_clk      => ad1939_subsystem_audio_fabric_system_clk_clk,        --    ad1939_subsystem_audio_fabric_system_clk.clk
			clk_reset_inputs_hps_clk_out_clk                  => clk_reset_inputs_hps_clk_out_clk,                    --                clk_reset_inputs_hps_clk_out.clk
			audio_mini_leds_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                  -- audio_mini_leds_reset_reset_bridge_in_reset.reset
			jtag_master_clk_reset_reset_bridge_in_reset_reset => rst_controller_003_reset_out_reset,                  -- jtag_master_clk_reset_reset_bridge_in_reset.reset
			Pitch_Shift_0_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                      --   Pitch_Shift_0_reset_reset_bridge_in_reset.reset
			system_id_reset_reset_bridge_in_reset_reset       => rst_controller_003_reset_out_reset,                  --       system_id_reset_reset_bridge_in_reset.reset
			jtag_master_master_address                        => jtag_master_master_address,                          --                          jtag_master_master.address
			jtag_master_master_waitrequest                    => jtag_master_master_waitrequest,                      --                                            .waitrequest
			jtag_master_master_byteenable                     => jtag_master_master_byteenable,                       --                                            .byteenable
			jtag_master_master_read                           => jtag_master_master_read,                             --                                            .read
			jtag_master_master_readdata                       => jtag_master_master_readdata,                         --                                            .readdata
			jtag_master_master_readdatavalid                  => jtag_master_master_readdatavalid,                    --                                            .readdatavalid
			jtag_master_master_write                          => jtag_master_master_write,                            --                                            .write
			jtag_master_master_writedata                      => jtag_master_master_writedata,                        --                                            .writedata
			audio_mini_leds_s1_address                        => mm_interconnect_0_audio_mini_leds_s1_address,        --                          audio_mini_leds_s1.address
			audio_mini_leds_s1_write                          => mm_interconnect_0_audio_mini_leds_s1_write,          --                                            .write
			audio_mini_leds_s1_readdata                       => mm_interconnect_0_audio_mini_leds_s1_readdata,       --                                            .readdata
			audio_mini_leds_s1_writedata                      => mm_interconnect_0_audio_mini_leds_s1_writedata,      --                                            .writedata
			audio_mini_leds_s1_chipselect                     => mm_interconnect_0_audio_mini_leds_s1_chipselect,     --                                            .chipselect
			de10_leds_s1_address                              => mm_interconnect_0_de10_leds_s1_address,              --                                de10_leds_s1.address
			de10_leds_s1_write                                => mm_interconnect_0_de10_leds_s1_write,                --                                            .write
			de10_leds_s1_readdata                             => mm_interconnect_0_de10_leds_s1_readdata,             --                                            .readdata
			de10_leds_s1_writedata                            => mm_interconnect_0_de10_leds_s1_writedata,            --                                            .writedata
			de10_leds_s1_chipselect                           => mm_interconnect_0_de10_leds_s1_chipselect,           --                                            .chipselect
			Pitch_Shift_0_avalon_mm_address                   => mm_interconnect_0_pitch_shift_0_avalon_mm_address,   --                     Pitch_Shift_0_avalon_mm.address
			Pitch_Shift_0_avalon_mm_write                     => mm_interconnect_0_pitch_shift_0_avalon_mm_write,     --                                            .write
			Pitch_Shift_0_avalon_mm_read                      => mm_interconnect_0_pitch_shift_0_avalon_mm_read,      --                                            .read
			Pitch_Shift_0_avalon_mm_readdata                  => mm_interconnect_0_pitch_shift_0_avalon_mm_readdata,  --                                            .readdata
			Pitch_Shift_0_avalon_mm_writedata                 => mm_interconnect_0_pitch_shift_0_avalon_mm_writedata, --                                            .writedata
			system_id_control_slave_address                   => mm_interconnect_0_system_id_control_slave_address,   --                     system_id_control_slave.address
			system_id_control_slave_readdata                  => mm_interconnect_0_system_id_control_slave_readdata   --                                            .readdata
		);

	rst_controller : component soc_system_passthrough_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => clk_reset_inputs_fabric_reset_out_reset,         -- reset_in0.reset
			reset_in1      => clk_reset_inputs_hps_and_fabric_reset_out_reset, -- reset_in1.reset
			clk            => ad1939_subsystem_audio_fabric_system_clk_clk,    --       clk.clk
			reset_out      => rst_controller_reset_out_reset,                  -- reset_out.reset
			reset_req      => open,                                            -- (terminated)
			reset_req_in0  => '0',                                             -- (terminated)
			reset_req_in1  => '0',                                             -- (terminated)
			reset_in2      => '0',                                             -- (terminated)
			reset_req_in2  => '0',                                             -- (terminated)
			reset_in3      => '0',                                             -- (terminated)
			reset_req_in3  => '0',                                             -- (terminated)
			reset_in4      => '0',                                             -- (terminated)
			reset_req_in4  => '0',                                             -- (terminated)
			reset_in5      => '0',                                             -- (terminated)
			reset_req_in5  => '0',                                             -- (terminated)
			reset_in6      => '0',                                             -- (terminated)
			reset_req_in6  => '0',                                             -- (terminated)
			reset_in7      => '0',                                             -- (terminated)
			reset_req_in7  => '0',                                             -- (terminated)
			reset_in8      => '0',                                             -- (terminated)
			reset_req_in8  => '0',                                             -- (terminated)
			reset_in9      => '0',                                             -- (terminated)
			reset_req_in9  => '0',                                             -- (terminated)
			reset_in10     => '0',                                             -- (terminated)
			reset_req_in10 => '0',                                             -- (terminated)
			reset_in11     => '0',                                             -- (terminated)
			reset_req_in11 => '0',                                             -- (terminated)
			reset_in12     => '0',                                             -- (terminated)
			reset_req_in12 => '0',                                             -- (terminated)
			reset_in13     => '0',                                             -- (terminated)
			reset_req_in13 => '0',                                             -- (terminated)
			reset_in14     => '0',                                             -- (terminated)
			reset_req_in14 => '0',                                             -- (terminated)
			reset_in15     => '0',                                             -- (terminated)
			reset_req_in15 => '0'                                              -- (terminated)
		);

	rst_controller_001 : component soc_system_passthrough_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => clk_reset_inputs_fabric_reset_out_reset,         -- reset_in0.reset
			reset_in1      => clk_reset_inputs_hps_and_fabric_reset_out_reset, -- reset_in1.reset
			clk            => open,                                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,              -- reset_out.reset
			reset_req      => open,                                            -- (terminated)
			reset_req_in0  => '0',                                             -- (terminated)
			reset_req_in1  => '0',                                             -- (terminated)
			reset_in2      => '0',                                             -- (terminated)
			reset_req_in2  => '0',                                             -- (terminated)
			reset_in3      => '0',                                             -- (terminated)
			reset_req_in3  => '0',                                             -- (terminated)
			reset_in4      => '0',                                             -- (terminated)
			reset_req_in4  => '0',                                             -- (terminated)
			reset_in5      => '0',                                             -- (terminated)
			reset_req_in5  => '0',                                             -- (terminated)
			reset_in6      => '0',                                             -- (terminated)
			reset_req_in6  => '0',                                             -- (terminated)
			reset_in7      => '0',                                             -- (terminated)
			reset_req_in7  => '0',                                             -- (terminated)
			reset_in8      => '0',                                             -- (terminated)
			reset_req_in8  => '0',                                             -- (terminated)
			reset_in9      => '0',                                             -- (terminated)
			reset_req_in9  => '0',                                             -- (terminated)
			reset_in10     => '0',                                             -- (terminated)
			reset_req_in10 => '0',                                             -- (terminated)
			reset_in11     => '0',                                             -- (terminated)
			reset_req_in11 => '0',                                             -- (terminated)
			reset_in12     => '0',                                             -- (terminated)
			reset_req_in12 => '0',                                             -- (terminated)
			reset_in13     => '0',                                             -- (terminated)
			reset_req_in13 => '0',                                             -- (terminated)
			reset_in14     => '0',                                             -- (terminated)
			reset_req_in14 => '0',                                             -- (terminated)
			reset_in15     => '0',                                             -- (terminated)
			reset_req_in15 => '0'                                              -- (terminated)
		);

	rst_controller_002 : component soc_system_passthrough_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => clk_reset_inputs_hps_and_fabric_reset_out_reset, -- reset_in0.reset
			clk            => clk_reset_inputs_hps_clk_out_clk,                --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,              -- reset_out.reset
			reset_req      => open,                                            -- (terminated)
			reset_req_in0  => '0',                                             -- (terminated)
			reset_in1      => '0',                                             -- (terminated)
			reset_req_in1  => '0',                                             -- (terminated)
			reset_in2      => '0',                                             -- (terminated)
			reset_req_in2  => '0',                                             -- (terminated)
			reset_in3      => '0',                                             -- (terminated)
			reset_req_in3  => '0',                                             -- (terminated)
			reset_in4      => '0',                                             -- (terminated)
			reset_req_in4  => '0',                                             -- (terminated)
			reset_in5      => '0',                                             -- (terminated)
			reset_req_in5  => '0',                                             -- (terminated)
			reset_in6      => '0',                                             -- (terminated)
			reset_req_in6  => '0',                                             -- (terminated)
			reset_in7      => '0',                                             -- (terminated)
			reset_req_in7  => '0',                                             -- (terminated)
			reset_in8      => '0',                                             -- (terminated)
			reset_req_in8  => '0',                                             -- (terminated)
			reset_in9      => '0',                                             -- (terminated)
			reset_req_in9  => '0',                                             -- (terminated)
			reset_in10     => '0',                                             -- (terminated)
			reset_req_in10 => '0',                                             -- (terminated)
			reset_in11     => '0',                                             -- (terminated)
			reset_req_in11 => '0',                                             -- (terminated)
			reset_in12     => '0',                                             -- (terminated)
			reset_req_in12 => '0',                                             -- (terminated)
			reset_in13     => '0',                                             -- (terminated)
			reset_req_in13 => '0',                                             -- (terminated)
			reset_in14     => '0',                                             -- (terminated)
			reset_req_in14 => '0',                                             -- (terminated)
			reset_in15     => '0',                                             -- (terminated)
			reset_req_in15 => '0'                                              -- (terminated)
		);

	rst_controller_003 : component soc_system_passthrough_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_h2f_reset_reset_ports_inv,      -- reset_in0.reset
			clk            => clk_reset_inputs_hps_clk_out_clk,   --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	hps_h2f_reset_reset_ports_inv <= not hps_h2f_reset_reset;

	clk_reset_inputs_hps_and_fabric_reset_out_reset_ports_inv <= not clk_reset_inputs_hps_and_fabric_reset_out_reset;

	mm_interconnect_0_audio_mini_leds_s1_write_ports_inv <= not mm_interconnect_0_audio_mini_leds_s1_write;

	mm_interconnect_0_de10_leds_s1_write_ports_inv <= not mm_interconnect_0_de10_leds_s1_write;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	rst_controller_003_reset_out_reset_ports_inv <= not rst_controller_003_reset_out_reset;

end architecture rtl; -- of soc_system_passthrough
