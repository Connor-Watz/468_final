-- soc_system_passthrough_clk_reset_inputs.vhd

-- Generated using ACDS version 21.1 842

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system_passthrough_clk_reset_inputs is
	port (
		fabric_reset_in_reset          : in  std_logic := '0'; --          fabric_reset_in.reset
		fabric_reset_out_reset         : out std_logic;        --         fabric_reset_out.reset
		hps_and_fabric_reset_in_reset  : in  std_logic := '0'; --  hps_and_fabric_reset_in.reset
		hps_and_fabric_reset_out_reset : out std_logic;        -- hps_and_fabric_reset_out.reset
		hps_clk_in_clk                 : in  std_logic := '0'; --               hps_clk_in.clk
		hps_clk_out_clk                : out std_logic         --              hps_clk_out.clk
	);
end entity soc_system_passthrough_clk_reset_inputs;

architecture rtl of soc_system_passthrough_clk_reset_inputs is
begin

	fabric_reset_out_reset <= fabric_reset_in_reset;

	hps_and_fabric_reset_out_reset <= hps_and_fabric_reset_in_reset;

	hps_clk_out_clk <= hps_clk_in_clk;

end architecture rtl; -- of soc_system_passthrough_clk_reset_inputs
